module extensor16para32(a, x);
input [15:0]a;
output [31:0]x;
assign x[0] = a[0];
assign x[1] = a[1];
assign x[2] = a[2];
assign x[3] = a[3];
assign x[4] = a[4];
assign x[5] = a[5];
assign x[6] = a[6];
assign x[7] = a[7];
assign x[8] = a[8];
assign x[9] = a[9];
assign x[10] = a[10];
assign x[11] = a[11];
assign x[12] = a[12];
assign x[13] = a[13];
assign x[14] = a[14];
assign x[15] = a[15];
assign x[16] = a[15];
assign x[17] = a[15];
assign x[18] = a[15];
assign x[19] = a[15];
assign x[20] = a[15];
assign x[21] = a[15];
assign x[22] = a[15];
assign x[23] = a[15];
assign x[24] = a[15];
assign x[25] = a[15];
assign x[26] = a[15];
assign x[27] = a[15];
assign x[28] = a[15];
assign x[29] = a[15];
assign x[30] = a[15];
assign x[31] = a[15];
endmodule