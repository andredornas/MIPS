library verilog;
use verilog.vl_types.all;
entity slt is
    port(
        a               : in     vl_logic_vector(31 downto 0);
        b               : in     vl_logic_vector(31 downto 0);
        x               : out    vl_logic_vector(31 downto 0)
    );
end slt;
